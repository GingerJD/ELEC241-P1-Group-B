module servo_control_unit_tb;

//Set initial variables for servo_control_unit.sv
logic Direction;
logic brake;
logic resetOut;
logic [7:0] pwmDT;
logic [7:0] pwmPeriod;
logic [31:0] statusR;
logic [31:0] inputR;
logic [11:0] atuAngle;

//Initialize servo_control_unit.sv

scu u1(Direction, brake, resetOut, pwmDT,pwmPeriod,statusR,inputR,atuAngle);
initial begin
inputR = 32'b10000000000011001000000000011100;
atuAngle = 576;	

#300 atuAngle = 12'b000000011100;
//////////////////////////////////////////////////////////////////////////////
//TEST 1 - Possile to set desired angle

//////////////////////////////////////////////////////////////////////////////
//TEST 2 - Bang Bang control

//////////////////////////////////////////////////////////////////////////////
//TEST 3 - Proortional control

//////////////////////////////////////////////////////////////////////////////
//TEST 4 - inputR is read correctly

//////////////////////////////////////////////////////////////////////////////
//TEST 5 - statusR is written correctly

//////////////////////////////////////////////////////////////////////////////
//TEST 6 - Current angle is output for DC 

//////////////////////////////////////////////////////////////////////////////
//TEST 7 - CONTINUOUS COMMAND TEST

//////////////////////////////////////////////////////////////////////////////
//TEST 8 - RESET COMMAND TEST

//////////////////////////////////////////////////////////////////////////////
//TEST 9 - NC COMMAND TEST

//////////////////////////////////////////////////////////////////////////////
//TEST 10 - BRAKE COMMAND TEST - NEEDS TO OVERRIDE PWM POWER











end
endmodule


